-- ========================================
-- [] File Name : network.vhdl
--
-- [] Creation Date : January 2018
--
-- [] Author 1 : Ali Gholami (aligholami7596@gmail.com)
--
-- [] Author 2 : Mehdi Safaee(mxii1994@gmail.com)
-- ========================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity BitonicSort is
    generic(NETWORK_BUS_WIDTH: INTEGER := 16);
    port(
        NET_INPUT: in 
    );
end BitonicSort;

architecture RTL of BitonicSort is

begin

end RTL;
